module sigmoid_lut (
    input clk,
    input reset,
    input signed [7:0] x_in,  // Q3.5 input (-4 to 4)
    output reg [7:0] y_out    // Q0.8 output (0 to 1)
);

     reg [7:0] LUT [255:0];

    //registering output
    always @(posedge clk or negedge reset) begin
      if(~reset) begin
        y_out <= 0;
      end
      else begin
        y_out <= LUT['sd128+x_in];
      end
    end 


    always @(posedge clk or negedge reset) begin
      LUT[0]  <= 5; LUT[1]  <= 5; LUT[2]  <= 5; LUT[3]  <= 5; LUT[4]  <= 5; LUT[5]  <= 5;
      LUT[6]  <= 6; LUT[7]  <= 6; LUT[8]  <= 6; LUT[9]  <= 6; LUT[10] <= 6; LUT[11] <= 6;
      LUT[12] <= 7; LUT[13] <= 7; LUT[14] <= 7; LUT[15] <= 7; LUT[16] <= 8; LUT[17] <= 8;
      LUT[18] <= 8; LUT[19] <= 8; LUT[20] <= 8; LUT[21] <= 9; LUT[22] <= 9; LUT[23] <= 9;
      LUT[24] <= 10; LUT[25] <= 10; LUT[26] <= 10; LUT[27] <= 10; LUT[28] <= 11; LUT[29] <= 11;
      LUT[30] <= 11; LUT[31] <= 12; LUT[32] <= 12; LUT[33] <= 13; LUT[34] <= 13; LUT[35] <= 13;
      LUT[36] <= 14; LUT[37] <= 14; LUT[38] <= 15; LUT[39] <= 15; LUT[40] <= 15; LUT[41] <= 16;
      LUT[42] <= 16; LUT[43] <= 17; LUT[44] <= 17; LUT[45] <= 18; LUT[46] <= 18; LUT[47] <= 19;
      LUT[48] <= 19; LUT[49] <= 20; LUT[50] <= 21; LUT[51] <= 21; LUT[52] <= 22; LUT[53] <= 22;
      LUT[54] <= 23; LUT[55] <= 24; LUT[56] <= 24; LUT[57] <= 25; LUT[58] <= 26; LUT[59] <= 27;
      LUT[60] <= 27; LUT[61] <= 28; LUT[62] <= 29; LUT[63] <= 30; LUT[64] <= 31; LUT[65] <= 31;
      LUT[66] <= 32; LUT[67] <= 33; LUT[68] <= 34; LUT[69] <= 35; LUT[70] <= 36; LUT[71] <= 37;
      LUT[72] <= 38; LUT[73] <= 39; LUT[74] <= 40; LUT[75] <= 41; LUT[76] <= 42; LUT[77] <= 43;
      LUT[78] <= 44; LUT[79] <= 46; LUT[80] <= 47; LUT[81] <= 48; LUT[82] <= 49; LUT[83] <= 50;
      LUT[84] <= 52; LUT[85] <= 53; LUT[86] <= 54; LUT[87] <= 56; LUT[88] <= 57; LUT[89] <= 58;
      LUT[90] <= 60; LUT[91] <= 61; LUT[92] <= 63; LUT[93] <= 64; LUT[94] <= 66; LUT[95] <= 67;
      LUT[96] <= 69; LUT[97] <= 70; LUT[98] <= 72; LUT[99] <= 74; LUT[100] <= 75; LUT[101] <= 77;
      LUT[102] <= 79; LUT[103] <= 80; LUT[104] <= 82; LUT[105] <= 84; LUT[106] <= 86; LUT[107] <= 87;
      LUT[108] <= 89; LUT[109] <= 91; LUT[110] <= 93; LUT[111] <= 95; LUT[112] <= 97; LUT[113] <= 99;
      LUT[114] <= 100; LUT[115] <= 102; LUT[116] <= 104; LUT[117] <= 106; LUT[118] <= 108; LUT[119] <= 110;
      LUT[120] <= 112; LUT[121] <= 114; LUT[122] <= 116; LUT[123] <= 118; LUT[124] <= 120; LUT[125] <= 122;
      LUT[126] <= 124; LUT[127] <= 126; LUT[128] <= 128; LUT[129] <= 130; LUT[130] <= 132; LUT[131] <= 134;
      LUT[132] <= 136; LUT[133] <= 138; LUT[134] <= 140; LUT[135] <= 142; LUT[136] <= 144; LUT[137] <= 146;
      LUT[138] <= 148; LUT[139] <= 150; LUT[140] <= 152; LUT[141] <= 154; LUT[142] <= 156; LUT[143] <= 157;
      LUT[144] <= 159; LUT[145] <= 161; LUT[146] <= 163; LUT[147] <= 165; LUT[148] <= 167; LUT[149] <= 169;
      LUT[150] <= 170; LUT[151] <= 172; LUT[152] <= 174; LUT[153] <= 176; LUT[154] <= 177; LUT[155] <= 179;
      LUT[156] <= 181; LUT[157] <= 182; LUT[158] <= 184; LUT[159] <= 186; LUT[160] <= 187; LUT[161] <= 189;
      LUT[162] <= 190; LUT[163] <= 192; LUT[164] <= 193; LUT[165] <= 195; LUT[166] <= 196; LUT[167] <= 198;
      LUT[168] <= 199; LUT[169] <= 200; LUT[170] <= 202; LUT[171] <= 203; LUT[172] <= 204; LUT[173] <= 206;
      LUT[174] <= 207; LUT[175] <= 208; LUT[176] <= 209; LUT[177] <= 210; LUT[178] <= 212; LUT[179] <= 213;
      LUT[180] <= 214; LUT[181] <= 215; LUT[182] <= 216; LUT[183] <= 217; LUT[184] <= 218; LUT[185] <= 219;
      LUT[186] <= 220; LUT[187] <= 221; LUT[188] <= 222; LUT[189] <= 223; LUT[190] <= 224; LUT[191] <= 225;
      LUT[192] <= 225; LUT[193] <= 226; LUT[194] <= 227; LUT[195] <= 228; LUT[196] <= 229; LUT[197] <= 229;
      LUT[198] <= 230; LUT[199] <= 231; LUT[200] <= 232; LUT[201] <= 232; LUT[202] <= 233; LUT[203] <= 234;
      LUT[204] <= 234; LUT[205] <= 235; LUT[206] <= 235; LUT[207] <= 236; LUT[208] <= 237; LUT[209] <= 237;
      LUT[210] <= 238; LUT[211] <= 238; LUT[212] <= 239; LUT[213] <= 239; LUT[214] <= 240; LUT[215] <= 240;
      LUT[216] <= 241; LUT[217] <= 241; LUT[218] <= 241; LUT[219] <= 242; LUT[220] <= 242; LUT[221] <= 243;
      LUT[222] <= 243; LUT[223] <= 243; LUT[224] <= 244; LUT[225] <= 244; LUT[226] <= 245; LUT[227] <= 245;
      LUT[228] <= 245; LUT[229] <= 246; LUT[230] <= 246; LUT[231] <= 246; LUT[232] <= 246; LUT[233] <= 247;
      LUT[234] <= 247; LUT[235] <= 247; LUT[236] <= 248; LUT[237] <= 248; LUT[238] <= 248; LUT[239] <= 248;
      LUT[240] <= 248; LUT[241] <= 249; LUT[242] <= 249; LUT[243] <= 249; LUT[244] <= 250; LUT[245] <= 250;
      LUT[246] <= 250; LUT[247] <= 250; LUT[248] <= 250; LUT[249] <= 250; LUT[250] <= 251; LUT[251] <= 251;
      LUT[252] <= 251; LUT[253] <= 251; LUT[254] <= 251; LUT[255] <= 251;
    end

endmodule

