module tanh_lut (
    input clk,
    input reset,
    input signed [7:0] x_in,  // Q3.5 input (-4 to 4)
    output reg signed [7:0] y_out    // Q0.7 output (-1 to 1)
);

     reg signed [7:0] LUT [255:0];

    //registering output
    always @(posedge clk or negedge reset) begin
      if(~reset) begin
        y_out <= 0;
      end
      else begin
        y_out <= LUT['sd128+x_in];
      end
    end 


    always @(posedge clk or negedge reset) begin
      LUT[0] <= -128;
      LUT[1] <= -128;
      LUT[2] <= -128;
      LUT[3] <= -128;
      LUT[4] <= -128;
      LUT[5] <= -128;
      LUT[6] <= -128;
      LUT[7] <= -128;
      LUT[8] <= -128;
      LUT[9] <= -128;
      LUT[10] <= -128;
      LUT[11] <= -128;
      LUT[12] <= -128;
      LUT[13] <= -128;
      LUT[14] <= -128;
      LUT[15] <= -128;
      LUT[16] <= -128;
      LUT[17] <= -128;
      LUT[18] <= -128;
      LUT[19] <= -128;
      LUT[20] <= -128;
      LUT[21] <= -128;
      LUT[22] <= -128;
      LUT[23] <= -128;
      LUT[24] <= -128;
      LUT[25] <= -128;
      LUT[26] <= -128;
      LUT[27] <= -128;
      LUT[28] <= -128;
      LUT[29] <= -127;
      LUT[30] <= -127;
      LUT[31] <= -127;
      LUT[32] <= -127;
      LUT[33] <= -127;
      LUT[34] <= -127;
      LUT[35] <= -127;
      LUT[36] <= -127;
      LUT[37] <= -127;
      LUT[38] <= -127;
      LUT[39] <= -127;
      LUT[40] <= -127;
      LUT[41] <= -127;
      LUT[42] <= -127;
      LUT[43] <= -127;
      LUT[44] <= -127;
      LUT[45] <= -126;
      LUT[46] <= -126;
      LUT[47] <= -126;
      LUT[48] <= -126;
      LUT[49] <= -126;
      LUT[50] <= -126;
      LUT[51] <= -126;
      LUT[52] <= -126;
      LUT[53] <= -126;
      LUT[54] <= -125;
      LUT[55] <= -125;
      LUT[56] <= -125;
      LUT[57] <= -125;
      LUT[58] <= -125;
      LUT[59] <= -124;
      LUT[60] <= -124;
      LUT[61] <= -124;
      LUT[62] <= -124;
      LUT[63] <= -123;
      LUT[64] <= -123;
      LUT[65] <= -123;
      LUT[66] <= -122;
      LUT[67] <= -122;
      LUT[68] <= -122;
      LUT[69] <= -121;
      LUT[70] <= -121;
      LUT[71] <= -120;
      LUT[72] <= -120;
      LUT[73] <= -120;
      LUT[74] <= -119;
      LUT[75] <= -118;
      LUT[76] <= -118;
      LUT[77] <= -117;
      LUT[78] <= -117;
      LUT[79] <= -116;
      LUT[80] <= -115;
      LUT[81] <= -114;
      LUT[82] <= -113;
      LUT[83] <= -113;
      LUT[84] <= -112;
      LUT[85] <= -111;
      LUT[86] <= -110;
      LUT[87] <= -109;
      LUT[88] <= -107;
      LUT[89] <= -106;
      LUT[90] <= -105;
      LUT[91] <= -104;
      LUT[92] <= -102;
      LUT[93] <= -101;
      LUT[94] <= -99;
      LUT[95] <= -97;
      LUT[96] <= -96;
      LUT[97] <= -94;
      LUT[98] <= -92;
      LUT[99] <= -90;
      LUT[100] <= -88;
      LUT[101] <= -86;
      LUT[102] <= -84;
      LUT[103] <= -81;
      LUT[104] <= -79;
      LUT[105] <= -76;
      LUT[106] <= -74;
      LUT[107] <= -71;
      LUT[108] <= -68;
      LUT[109] <= -65;
      LUT[110] <= -62;
      LUT[111] <= -59;
      LUT[112] <= -56;
      LUT[113] <= -53;
      LUT[114] <= -49;
      LUT[115] <= -46;
      LUT[116] <= -42;
      LUT[117] <= -39;
      LUT[118] <= -35;
      LUT[119] <= -31;
      LUT[120] <= -28;
      LUT[121] <= -24;
      LUT[122] <= -20;
      LUT[123] <= -16;
      LUT[124] <= -12;
      LUT[125] <= -8;
      LUT[126] <= -4;
      LUT[127] <= 0;
      LUT[128] <= 4;
      LUT[129] <= 8;
      LUT[130] <= 12;
      LUT[131] <= 16;
      LUT[132] <= 20;
      LUT[133] <= 24;
      LUT[134] <= 28;
      LUT[135] <= 31;
      LUT[136] <= 35;
      LUT[137] <= 39;
      LUT[138] <= 42;
      LUT[139] <= 46;
      LUT[140] <= 49;
      LUT[141] <= 53;
      LUT[142] <= 56;
      LUT[143] <= 59;
      LUT[144] <= 62;
      LUT[145] <= 65;
      LUT[146] <= 68;
      LUT[147] <= 71;
      LUT[148] <= 74;
      LUT[149] <= 76;
      LUT[150] <= 79;
      LUT[151] <= 81;
      LUT[152] <= 84;
      LUT[153] <= 86;
      LUT[154] <= 88;
      LUT[155] <= 90;
      LUT[156] <= 92;
      LUT[157] <= 94;
      LUT[158] <= 96;
      LUT[159] <= 97;
      LUT[160] <= 99;
      LUT[161] <= 101;
      LUT[162] <= 102;
      LUT[163] <= 104;
      LUT[164] <= 105;
      LUT[165] <= 106;
      LUT[166] <= 107;
      LUT[167] <= 109;
      LUT[168] <= 110;
      LUT[169] <= 111;
      LUT[170] <= 112;
      LUT[171] <= 113;
      LUT[172] <= 113;
      LUT[173] <= 114;
      LUT[174] <= 115;
      LUT[175] <= 116;
      LUT[176] <= 117;
      LUT[177] <= 117;
      LUT[178] <= 118;
      LUT[179] <= 118;
      LUT[180] <= 119;
      LUT[181] <= 120;
      LUT[182] <= 120;
      LUT[183] <= 120;
      LUT[184] <= 121;
      LUT[185] <= 121;
      LUT[186] <= 122;
      LUT[187] <= 122;
      LUT[188] <= 122;
      LUT[189] <= 123;
      LUT[190] <= 123;
      LUT[191] <= 123;
      LUT[192] <= 124;
      LUT[193] <= 124;
      LUT[194] <= 124;
      LUT[195] <= 124;
      LUT[196] <= 125;
      LUT[197] <= 125;
      LUT[198] <= 125;
      LUT[199] <= 125;
      LUT[200] <= 125;
      LUT[201] <= 126;
      LUT[202] <= 126;
      LUT[203] <= 126;
      LUT[204] <= 126;
      LUT[205] <= 126;
      LUT[206] <= 126;
      LUT[207] <= 126;
      LUT[208] <= 126;
      LUT[209] <= 126;
      LUT[210] <= 127;
      LUT[211] <= 127;
      LUT[212] <= 127;
      LUT[213] <= 127;
      LUT[214] <= 127;
      LUT[215] <= 127;
      LUT[216] <= 127;
      LUT[217] <= 127;
      LUT[218] <= 127;
      LUT[219] <= 127;
      LUT[220] <= 127;
      LUT[221] <= 127;
      LUT[222] <= 127;
      LUT[223] <= 127;
      LUT[224] <= 127;
      LUT[225] <= 127;
      LUT[226] <= 127;
      LUT[227] <= 127;
      LUT[228] <= 127;
      LUT[229] <= 127;
      LUT[230] <= 127;
      LUT[231] <= 127;
      LUT[232] <= 127;
      LUT[233] <= 127;
      LUT[234] <= 127;
      LUT[235] <= 127;
      LUT[236] <= 127;
      LUT[237] <= 127;
      LUT[238] <= 127;
      LUT[239] <= 127;
      LUT[240] <= 127;
      LUT[241] <= 127;
      LUT[242] <= 127;
      LUT[243] <= 127;
      LUT[244] <= 127;
      LUT[245] <= 127;
      LUT[246] <= 127;
      LUT[247] <= 127;
      LUT[248] <= 127;
      LUT[249] <= 127;
      LUT[250] <= 127;
      LUT[251] <= 127;
      LUT[252] <= 127;
      LUT[253] <= 127;
      LUT[254] <= 127;
      LUT[255] <= 127;
    end

endmodule


