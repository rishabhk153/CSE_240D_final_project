module gelu_lut (
    input clk,
    input reset,
    input signed [7:0] x_in,  // Q3.5 input (-4 to 4)
    output reg signed [7:0] y_out    // Q3.5 output (-4 to 4)
);

     reg signed [7:0] LUT [255:0];

    //registering output
    always @(posedge clk or negedge reset) begin
      if(~reset) begin
        y_out <= 0;
      end
      else begin
        y_out <= LUT['sd128+x_in];
      end
    end 


    always @(posedge clk or negedge reset) begin
      LUT[0]<=0;
      LUT[1]<=0;
      LUT[2]<=0;
      LUT[3]<=0;
      LUT[4]<=0;
      LUT[5]<=0;
      LUT[6]<=0;
      LUT[7]<=0;
      LUT[8]<=0;
      LUT[9]<=0;
      LUT[10]<=0;
      LUT[11]<=0;
      LUT[12]<=0;
      LUT[13]<=0;
      LUT[14]<=0;
      LUT[15]<=0;
      LUT[16]<=0;
      LUT[17]<=0;
      LUT[18]<=0;
      LUT[19]<=0;
      LUT[20]<=0;
      LUT[21]<=0;
      LUT[22]<=0;
      LUT[23]<=0;
      LUT[24]<=0;
      LUT[25]<=0;
      LUT[26]<=0;
      LUT[27]<=0;
      LUT[28]<=0;
      LUT[29]<=0;
      LUT[30]<=0;
      LUT[31]<=0;
      LUT[32]<=0;
      LUT[33]<=0;
      LUT[34]<=0;
      LUT[35]<=0;
      LUT[36]<=0;
      LUT[37]<=0;
      LUT[38]<=0;
      LUT[39]<=0;
      LUT[40]<=0;
      LUT[41]<=0;
      LUT[42]<=0;
      LUT[43]<=0;
      LUT[44]<=0;
      LUT[45]<=0;
      LUT[46]<=0;
      LUT[47]<=0;
      LUT[48]<=0;
      LUT[49]<=-1;
      LUT[50]<=-1;
      LUT[51]<=-1;
      LUT[52]<=-1;
      LUT[53]<=-1;
      LUT[54]<=-1;
      LUT[55]<=-1;
      LUT[56]<=-1;
      LUT[57]<=-1;
      LUT[58]<=-1;
      LUT[59]<=-1;
      LUT[60]<=-1;
      LUT[61]<=-1;
      LUT[62]<=-1;
      LUT[63]<=-1;
      LUT[64]<=-1;
      LUT[65]<=-2;
      LUT[66]<=-2;
      LUT[67]<=-2;
      LUT[68]<=-2;
      LUT[69]<=-2;
      LUT[70]<=-2;
      LUT[71]<=-2;
      LUT[72]<=-2;
      LUT[73]<=-2;
      LUT[74]<=-2;
      LUT[75]<=-3;
      LUT[76]<=-3;
      LUT[77]<=-3;
      LUT[78]<=-3;
      LUT[79]<=-3;
      LUT[80]<=-3;
      LUT[81]<=-3;
      LUT[82]<=-3;
      LUT[83]<=-4;
      LUT[84]<=-4;
      LUT[85]<=-4;
      LUT[86]<=-4;
      LUT[87]<=-4;
      LUT[88]<=-4;
      LUT[89]<=-4;
      LUT[90]<=-4;
      LUT[91]<=-5;
      LUT[92]<=-5;
      LUT[93]<=-5;
      LUT[94]<=-5;
      LUT[95]<=-5;
      LUT[96]<=-5;
      LUT[97]<=-5;
      LUT[98]<=-5;
      LUT[99]<=-5;
      LUT[100]<=-5;
      LUT[101]<=-5;
      LUT[102]<=-5;
      LUT[103]<=-5;
      LUT[104]<=-5;
      LUT[105]<=-5;
      LUT[106]<=-5;
      LUT[107]<=-5;
      LUT[108]<=-5;
      LUT[109]<=-5;
      LUT[110]<=-5;
      LUT[111]<=-5;
      LUT[112]<=-5;
      LUT[113]<=-5;
      LUT[114]<=-5;
      LUT[115]<=-4;
      LUT[116]<=-4;
      LUT[117]<=-4;
      LUT[118]<=-4;
      LUT[119]<=-4;
      LUT[120]<=-3;
      LUT[121]<=-3;
      LUT[122]<=-3;
      LUT[123]<=-2;
      LUT[124]<=-2;
      LUT[125]<=-1;
      LUT[126]<=-1;
      LUT[127]<=0;
      LUT[128]<=0;
      LUT[129]<=1;
      LUT[130]<=1;
      LUT[131]<=2;
      LUT[132]<=2;
      LUT[133]<=3;
      LUT[134]<=3;
      LUT[135]<=4;
      LUT[136]<=5;
      LUT[137]<=5;
      LUT[138]<=6;
      LUT[139]<=7;
      LUT[140]<=8;
      LUT[141]<=9;
      LUT[142]<=9;
      LUT[143]<=10;
      LUT[144]<=11;
      LUT[145]<=12;
      LUT[146]<=13;
      LUT[147]<=14;
      LUT[148]<=15;
      LUT[149]<=16;
      LUT[150]<=17;
      LUT[151]<=18;
      LUT[152]<=19;
      LUT[153]<=20;
      LUT[154]<=21;
      LUT[155]<=22;
      LUT[156]<=23;
      LUT[157]<=24;
      LUT[158]<=25;
      LUT[159]<=26;
      LUT[160]<=27;
      LUT[161]<=28;
      LUT[162]<=29;
      LUT[163]<=30;
      LUT[164]<=31;
      LUT[165]<=32;
      LUT[166]<=34;
      LUT[167]<=35;
      LUT[168]<=36;
      LUT[169]<=37;
      LUT[170]<=38;
      LUT[171]<=39;
      LUT[172]<=40;
      LUT[173]<=41;
      LUT[174]<=43;
      LUT[175]<=44;
      LUT[176]<=45;
      LUT[177]<=46;
      LUT[178]<=47;
      LUT[179]<=48;
      LUT[180]<=49;
      LUT[181]<=50;
      LUT[182]<=52;
      LUT[183]<=53;
      LUT[184]<=54;
      LUT[185]<=55;
      LUT[186]<=56;
      LUT[187]<=57;
      LUT[188]<=58;
      LUT[189]<=59;
      LUT[190]<=60;
      LUT[191]<=61;
      LUT[192]<=63;
      LUT[193]<=64;
      LUT[194]<=65;
      LUT[195]<=66;
      LUT[196]<=67;
      LUT[197]<=68;
      LUT[198]<=69;
      LUT[199]<=70;
      LUT[200]<=71;
      LUT[201]<=72;
      LUT[202]<=73;
      LUT[203]<=74;
      LUT[204]<=75;
      LUT[205]<=76;
      LUT[206]<=77;
      LUT[207]<=78;
      LUT[208]<=80;
      LUT[209]<=81;
      LUT[210]<=82;
      LUT[211]<=83;
      LUT[212]<=84;
      LUT[213]<=85;
      LUT[214]<=86;
      LUT[215]<=87;
      LUT[216]<=88;
      LUT[217]<=89;
      LUT[218]<=90;
      LUT[219]<=91;
      LUT[220]<=92;
      LUT[221]<=93;
      LUT[222]<=94;
      LUT[223]<=95;
      LUT[224]<=96;
      LUT[225]<=97;
      LUT[226]<=98;
      LUT[227]<=99;
      LUT[228]<=100;
      LUT[229]<=101;
      LUT[230]<=102;
      LUT[231]<=103;
      LUT[232]<=104;
      LUT[233]<=105;
      LUT[234]<=106;
      LUT[235]<=107;
      LUT[236]<=108;
      LUT[237]<=109;
      LUT[238]<=110;
      LUT[239]<=111;
      LUT[240]<=112;
      LUT[241]<=113;
      LUT[242]<=114;
      LUT[243]<=115;
      LUT[244]<=116;
      LUT[245]<=117;
      LUT[246]<=118;
      LUT[247]<=119;
      LUT[248]<=120;
      LUT[249]<=121;
      LUT[250]<=122;
      LUT[251]<=123;
      LUT[252]<=124;
      LUT[253]<=125;
      LUT[254]<=126;
      LUT[255]<=127;
      LUT[255]<=127;
    end

endmodule


